package simpleadder_pkg;
	import uvm_pkg::*;
	`include "C:/Users/HP/WORK_UVM/uvm-1.2/src/uvm_macros.svh" // added this with full path  

	`include "C:/Users/HP/WORK_MODELSIM/project_uvm_adder/simpleadder_sequencer.sv"
	`include "C:/Users/HP/WORK_MODELSIM/project_uvm_adder/simpleadder_monitor.sv"
	`include "C:/Users/HP/WORK_MODELSIM/project_uvm_adder/simpleadder_driver.sv"
	`include "C:/Users/HP/WORK_MODELSIM/project_uvm_adder/simpleadder_agent.sv"
	`include "C:/Users/HP/WORK_MODELSIM/project_uvm_adder/simpleadder_scoreboard.sv"
	`include "C:/Users/HP/WORK_MODELSIM/project_uvm_adder/simpleadder_config.sv"
	`include "C:/Users/HP/WORK_MODELSIM/project_uvm_adder/simpleadder_env.sv"
	`include "C:/Users/HP/WORK_MODELSIM/project_uvm_adder/simpleadder_test.sv"
endpackage: simpleadder_pkg